module tb_or_gate(
    reg a, b
    output wire y
);

endmodule